* Test netlist 1 -- appears in Lecture on static element stamps

R1 1 0 5
G2 1 0 1 2 2
C3 1 2 6
R4 2 0 8
Is 0 2 10

.end
